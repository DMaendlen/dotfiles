Vim�UnDo� �N,l�� �A���� Wh[�c��9�8�f�,��C   �                                   S��z    _�                     �        ����                                                                                                                                                                                                                                                                                                                                                             S��x     �   �   �               5�_�                    �        ����                                                                                                                                                                                                                                                                                                                                                             S��x     �   �   �               5�_�                     �        ����                                                                                                                                                                                                                                                                                                                                                             S��y    �   �   �           5��